--> Refer to Instruction register
